library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

use std.textio.all;
use ieee.std_logic_textio.all;

entity rom_eight_bit_magnitude_adder is
   Generic(
        DATA_WIDTH : integer:=8;
        ADDR_WIDTH : integer:=16
   );
   Port ( clk : in STD_LOGIC;
          a : in STD_LOGIC_VECTOR (DATA_WIDTH-1 downto 0);
          b : in STD_LOGIC_VECTOR (DATA_WIDTH-1 downto 0);
          sum : out STD_LOGIC_VECTOR (DATA_WIDTH downto 0));
end rom_eight_bit_magnitude_adder;

architecture Behavioral of rom_eight_bit_magnitude_adder is

constant ROM_DEPTH : integer := 2**ADDR_WIDTH;
type rom_type is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH downto 0);

    impure function init_rom return rom_type is
        file text_file_16_bit : text open READ_MODE is "sixteen-bit-rom.txt";
        variable text_line : line;
        variable rom_content : rom_type ;
        variable value: std_logic_vector(DATA_WIDTH downto 0);

        begin

            for i in 0 to ROM_DEPTH -1 loop
                readline(text_file_16_bit, text_line);
                read(text_line, value);
                rom_content(i) := value;
            end loop;
        return rom_content;
    end function;

signal addr_r : STD_LOGIC_VECTOR ((DATA_WIDTH * 2) - 1 downto 0);
signal rom_file: rom_type := init_rom;
signal rom: rom_type := (
    "000000000",
"000000001",
"000000010",
"000000011",
"000000100",
"000000101",
"000000110",
"000000111",
"000001000",
"000001001",
"000001010",
"000001011",
"000001100",
"000001101",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111110",
"101111111",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"101110010",
"001110011",
"101110100",
"001110101",
"101110110",
"001110111",
"101111000",
"001111001",
"101111010",
"001111011",
"101111100",
"001111101",
"101111110",
"001111111",
"000000001",
"000000010",
"000000011",
"000000100",
"000000101",
"000000110",
"000000111",
"000001000",
"000001001",
"000001010",
"000001011",
"000001100",
"000001101",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"110000000",
"110000000",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"101110001",
"001110010",
"101110011",
"001110100",
"101110101",
"001110110",
"101110111",
"001111000",
"101111001",
"001111010",
"101111011",
"001111100",
"101111101",
"001111110",
"000000010",
"000000011",
"000000100",
"000000101",
"000000110",
"000000111",
"000001000",
"000001001",
"000001010",
"000001011",
"000001100",
"000001101",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"101110010",
"001110011",
"101110100",
"001110101",
"101110110",
"001110111",
"101111000",
"001111001",
"101111010",
"001111011",
"101111100",
"001111101",
"000000011",
"000000100",
"000000101",
"000000110",
"000000111",
"000001000",
"000001001",
"000001010",
"000001011",
"000001100",
"000001101",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"110000010",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"101110001",
"001110010",
"101110011",
"001110100",
"101110101",
"001110110",
"101110111",
"001111000",
"101111001",
"001111010",
"101111011",
"001111100",
"000000100",
"000000101",
"000000110",
"000000111",
"000001000",
"000001001",
"000001010",
"000001011",
"000001100",
"000001101",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"101110010",
"001110011",
"101110100",
"001110101",
"101110110",
"001110111",
"101111000",
"001111001",
"101111010",
"001111011",
"000000101",
"000000110",
"000000111",
"000001000",
"000001001",
"000001010",
"000001011",
"000001100",
"000001101",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"110000100",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"101110001",
"001110010",
"101110011",
"001110100",
"101110101",
"001110110",
"101110111",
"001111000",
"101111001",
"001111010",
"000000110",
"000000111",
"000001000",
"000001001",
"000001010",
"000001011",
"000001100",
"000001101",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"101110010",
"001110011",
"101110100",
"001110101",
"101110110",
"001110111",
"101111000",
"001111001",
"000000111",
"000001000",
"000001001",
"000001010",
"000001011",
"000001100",
"000001101",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"110000110",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"101110001",
"001110010",
"101110011",
"001110100",
"101110101",
"001110110",
"101110111",
"001111000",
"000001000",
"000001001",
"000001010",
"000001011",
"000001100",
"000001101",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"101110010",
"001110011",
"101110100",
"001110101",
"101110110",
"001110111",
"000001001",
"000001010",
"000001011",
"000001100",
"000001101",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"110001000",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"101110001",
"001110010",
"101110011",
"001110100",
"101110101",
"001110110",
"000001010",
"000001011",
"000001100",
"000001101",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"101110010",
"001110011",
"101110100",
"001110101",
"000001011",
"000001100",
"000001101",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"110001010",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"101110001",
"001110010",
"101110011",
"001110100",
"000001100",
"000001101",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"101110010",
"001110011",
"000001101",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"110001100",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"101110001",
"001110010",
"000001110",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"000001111",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"110001110",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"000010000",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"000010001",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"110010000",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"000010010",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"000010011",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"110010010",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"000010100",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"000010101",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"110010100",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"000010110",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"000010111",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"110010110",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"000011000",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"000011001",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"110011000",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"000011010",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"000011011",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"110011010",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"000011100",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"000011101",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"110011100",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"000011110",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"000011111",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"110011110",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"000100000",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"000100001",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"110100000",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"000100010",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"000100011",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"110100010",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"000100100",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"000100101",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"110100100",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"000100110",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"000100111",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"110100110",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"000101000",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"000101001",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"110101000",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"000101010",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"000101011",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"110101010",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"000101100",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"000101101",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"110101100",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"000101110",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"000101111",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"110101110",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"000110000",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"000110001",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"110110000",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"000110010",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"000110011",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"110110010",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"000110100",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"000110101",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"110110100",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"000110110",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"000110111",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"110110110",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"000111000",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"000111001",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"110111000",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"000111010",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"000111011",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"110111010",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"000111100",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"000111101",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"110111100",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"000111110",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"000111111",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"110111110",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"001000000",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"001000001",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"111000000",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"001000010",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"001000011",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"111000010",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"001000100",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"001000101",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"111000100",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"001000110",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"001000111",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"111000110",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"001001000",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"001001001",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"111001000",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"001001010",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"001001011",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"111001010",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"001001100",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"001001101",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"111001100",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"001001110",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"001001111",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"111001110",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"001010000",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"001010001",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"111010000",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"001010010",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"001010011",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"111010010",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"001010100",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"001010101",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"111010100",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"001010110",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"001010111",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"111010110",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"001011000",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"001011001",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"111011000",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"001011010",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"001011011",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"111011010",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"001011100",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"001011101",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"111011100",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"001011110",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"001011111",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"111011110",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"001100000",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"001100001",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"111100000",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"001100010",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"001100011",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"111100010",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"001100100",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"001100101",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"111100100",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"001100110",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"001100111",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"111100110",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"001101000",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"001101001",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"111101000",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"001101010",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"001101011",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"111101010",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"001101100",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"001101101",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"111101100",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"001101110",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"001101111",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"111101110",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"001110000",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"001110001",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"111110000",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"001110010",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"011110000",
"011110001",
"001110010",
"001110001",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"001110011",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"011110000",
"011110001",
"111110010",
"101110011",
"101110010",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"001110100",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"011110000",
"011110001",
"011110010",
"011110011",
"001110100",
"001110011",
"001110010",
"001110001",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"001110101",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"011110000",
"011110001",
"011110010",
"011110011",
"111110100",
"101110101",
"101110100",
"101110011",
"101110010",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"001110110",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"011110000",
"011110001",
"011110010",
"011110011",
"011110100",
"011110101",
"001110110",
"001110101",
"001110100",
"001110011",
"001110010",
"001110001",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"001110111",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"011110000",
"011110001",
"011110010",
"011110011",
"011110100",
"011110101",
"111110110",
"101110111",
"101110110",
"101110101",
"101110100",
"101110011",
"101110010",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"001111000",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"011110000",
"011110001",
"011110010",
"011110011",
"011110100",
"011110101",
"011110110",
"011110111",
"001111000",
"001110111",
"001110110",
"001110101",
"001110100",
"001110011",
"001110010",
"001110001",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"001111001",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"011110000",
"011110001",
"011110010",
"011110011",
"011110100",
"011110101",
"011110110",
"011110111",
"111111000",
"101111001",
"101111000",
"101110111",
"101110110",
"101110101",
"101110100",
"101110011",
"101110010",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"001111010",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"011110000",
"011110001",
"011110010",
"011110011",
"011110100",
"011110101",
"011110110",
"011110111",
"011111000",
"011111001",
"001111010",
"001111001",
"001111000",
"001110111",
"001110110",
"001110101",
"001110100",
"001110011",
"001110010",
"001110001",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"001111011",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"011110000",
"011110001",
"011110010",
"011110011",
"011110100",
"011110101",
"011110110",
"011110111",
"011111000",
"011111001",
"111111010",
"101111011",
"101111010",
"101111001",
"101111000",
"101110111",
"101110110",
"101110101",
"101110100",
"101110011",
"101110010",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"001111100",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"011110000",
"011110001",
"011110010",
"011110011",
"011110100",
"011110101",
"011110110",
"011110111",
"011111000",
"011111001",
"011111010",
"011111011",
"001111100",
"001111011",
"001111010",
"001111001",
"001111000",
"001110111",
"001110110",
"001110101",
"001110100",
"001110011",
"001110010",
"001110001",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"001111101",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"011110000",
"011110001",
"011110010",
"011110011",
"011110100",
"011110101",
"011110110",
"011110111",
"011111000",
"011111001",
"011111010",
"011111011",
"111111100",
"101111101",
"101111100",
"101111011",
"101111010",
"101111001",
"101111000",
"101110111",
"101110110",
"101110101",
"101110100",
"101110011",
"101110010",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"001111110",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"011110000",
"011110001",
"011110010",
"011110011",
"011110100",
"011110101",
"011110110",
"011110111",
"011111000",
"011111001",
"011111010",
"011111011",
"011111100",
"011111101",
"001111110",
"001111101",
"001111100",
"001111011",
"001111010",
"001111001",
"001111000",
"001110111",
"001110110",
"001110101",
"001110100",
"001110011",
"001110010",
"001110001",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"001111111",
"010000000",
"010000001",
"010000010",
"010000011",
"010000100",
"010000101",
"010000110",
"010000111",
"010001000",
"010001001",
"010001010",
"010001011",
"010001100",
"010001101",
"010001110",
"010001111",
"010010000",
"010010001",
"010010010",
"010010011",
"010010100",
"010010101",
"010010110",
"010010111",
"010011000",
"010011001",
"010011010",
"010011011",
"010011100",
"010011101",
"010011110",
"010011111",
"010100000",
"010100001",
"010100010",
"010100011",
"010100100",
"010100101",
"010100110",
"010100111",
"010101000",
"010101001",
"010101010",
"010101011",
"010101100",
"010101101",
"010101110",
"010101111",
"010110000",
"010110001",
"010110010",
"010110011",
"010110100",
"010110101",
"010110110",
"010110111",
"010111000",
"010111001",
"010111010",
"010111011",
"010111100",
"010111101",
"010111110",
"010111111",
"011000000",
"011000001",
"011000010",
"011000011",
"011000100",
"011000101",
"011000110",
"011000111",
"011001000",
"011001001",
"011001010",
"011001011",
"011001100",
"011001101",
"011001110",
"011001111",
"011010000",
"011010001",
"011010010",
"011010011",
"011010100",
"011010101",
"011010110",
"011010111",
"011011000",
"011011001",
"011011010",
"011011011",
"011011100",
"011011101",
"011011110",
"011011111",
"011100000",
"011100001",
"011100010",
"011100011",
"011100100",
"011100101",
"011100110",
"011100111",
"011101000",
"011101001",
"011101010",
"011101011",
"011101100",
"011101101",
"011101110",
"011101111",
"011110000",
"011110001",
"011110010",
"011110011",
"011110100",
"011110101",
"011110110",
"011110111",
"011111000",
"011111001",
"011111010",
"011111011",
"011111100",
"011111101",
"111111110",
"101111111",
"101111110",
"101111101",
"101111100",
"101111011",
"101111010",
"101111001",
"101111000",
"101110111",
"101110110",
"101110101",
"101110100",
"101110011",
"101110010",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"100000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"101110010",
"001110011",
"101110100",
"001110101",
"101110110",
"001110111",
"101111000",
"001111001",
"101111010",
"001111011",
"101111100",
"001111101",
"101111110",
"101111111",
"100000000",
"100000001",
"100000010",
"100000011",
"100000100",
"100000101",
"100000110",
"100000111",
"100001000",
"100001001",
"100001010",
"100001011",
"100001100",
"100001101",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"101111111",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"101110001",
"001110010",
"101110011",
"001110100",
"101110101",
"001110110",
"101110111",
"001111000",
"101111001",
"001111010",
"101111011",
"001111100",
"101111101",
"101111110",
"100000001",
"100000010",
"100000011",
"100000100",
"100000101",
"100000110",
"100000111",
"100001000",
"100001001",
"100001010",
"100001011",
"100001100",
"100001101",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"010000000",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"101110010",
"001110011",
"101110100",
"001110101",
"101110110",
"001110111",
"101111000",
"001111001",
"101111010",
"001111011",
"101111100",
"101111101",
"100000010",
"100000011",
"100000100",
"100000101",
"100000110",
"100000111",
"100001000",
"100001001",
"100001010",
"100001011",
"100001100",
"100001101",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"101110001",
"001110010",
"101110011",
"001110100",
"101110101",
"001110110",
"101110111",
"001111000",
"101111001",
"001111010",
"101111011",
"101111100",
"100000011",
"100000100",
"100000101",
"100000110",
"100000111",
"100001000",
"100001001",
"100001010",
"100001011",
"100001100",
"100001101",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"010000010",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"101110010",
"001110011",
"101110100",
"001110101",
"101110110",
"001110111",
"101111000",
"001111001",
"101111010",
"101111011",
"100000100",
"100000101",
"100000110",
"100000111",
"100001000",
"100001001",
"100001010",
"100001011",
"100001100",
"100001101",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"101110001",
"001110010",
"101110011",
"001110100",
"101110101",
"001110110",
"101110111",
"001111000",
"101111001",
"101111010",
"100000101",
"100000110",
"100000111",
"100001000",
"100001001",
"100001010",
"100001011",
"100001100",
"100001101",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"010000100",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"101110010",
"001110011",
"101110100",
"001110101",
"101110110",
"001110111",
"101111000",
"101111001",
"100000110",
"100000111",
"100001000",
"100001001",
"100001010",
"100001011",
"100001100",
"100001101",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"101110001",
"001110010",
"101110011",
"001110100",
"101110101",
"001110110",
"101110111",
"101111000",
"100000111",
"100001000",
"100001001",
"100001010",
"100001011",
"100001100",
"100001101",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"010000110",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"101110010",
"001110011",
"101110100",
"001110101",
"101110110",
"101110111",
"100001000",
"100001001",
"100001010",
"100001011",
"100001100",
"100001101",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"101110001",
"001110010",
"101110011",
"001110100",
"101110101",
"101110110",
"100001001",
"100001010",
"100001011",
"100001100",
"100001101",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"010001000",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"101110010",
"001110011",
"101110100",
"101110101",
"100001010",
"100001011",
"100001100",
"100001101",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"101110001",
"001110010",
"101110011",
"101110100",
"100001011",
"100001100",
"100001101",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"010001010",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"001110001",
"101110010",
"101110011",
"100001100",
"100001101",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"001110000",
"101110001",
"101110010",
"100001101",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"010001100",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"001101111",
"101110000",
"101110001",
"100001110",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"001101110",
"101101111",
"101110000",
"100001111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"010001110",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"001101101",
"101101110",
"101101111",
"100010000",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"001101100",
"101101101",
"101101110",
"100010001",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"010010000",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"001101011",
"101101100",
"101101101",
"100010010",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"001101010",
"101101011",
"101101100",
"100010011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"010010010",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"001101001",
"101101010",
"101101011",
"100010100",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"001101000",
"101101001",
"101101010",
"100010101",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"010010100",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"001100111",
"101101000",
"101101001",
"100010110",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"001100110",
"101100111",
"101101000",
"100010111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"010010110",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"001100101",
"101100110",
"101100111",
"100011000",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"001100100",
"101100101",
"101100110",
"100011001",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"010011000",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"001100011",
"101100100",
"101100101",
"100011010",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"001100010",
"101100011",
"101100100",
"100011011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"010011010",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"001100001",
"101100010",
"101100011",
"100011100",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"001100000",
"101100001",
"101100010",
"100011101",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"010011100",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"001011111",
"101100000",
"101100001",
"100011110",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"001011110",
"101011111",
"101100000",
"100011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"010011110",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"001011101",
"101011110",
"101011111",
"100100000",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"001011100",
"101011101",
"101011110",
"100100001",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"010100000",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"001011011",
"101011100",
"101011101",
"100100010",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"001011010",
"101011011",
"101011100",
"100100011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"010100010",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"001011001",
"101011010",
"101011011",
"100100100",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"001011000",
"101011001",
"101011010",
"100100101",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"010100100",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"001010111",
"101011000",
"101011001",
"100100110",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"001010110",
"101010111",
"101011000",
"100100111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"010100110",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"001010101",
"101010110",
"101010111",
"100101000",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"001010100",
"101010101",
"101010110",
"100101001",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"010101000",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"001010011",
"101010100",
"101010101",
"100101010",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"001010010",
"101010011",
"101010100",
"100101011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"010101010",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"001010001",
"101010010",
"101010011",
"100101100",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"001010000",
"101010001",
"101010010",
"100101101",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"010101100",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"001001111",
"101010000",
"101010001",
"100101110",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"001001110",
"101001111",
"101010000",
"100101111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"010101110",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"001001101",
"101001110",
"101001111",
"100110000",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"001001100",
"101001101",
"101001110",
"100110001",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"010110000",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"001001011",
"101001100",
"101001101",
"100110010",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"001001010",
"101001011",
"101001100",
"100110011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"010110010",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"001001001",
"101001010",
"101001011",
"100110100",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"001001000",
"101001001",
"101001010",
"100110101",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"010110100",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"001000111",
"101001000",
"101001001",
"100110110",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"001000110",
"101000111",
"101001000",
"100110111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"010110110",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"001000101",
"101000110",
"101000111",
"100111000",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"001000100",
"101000101",
"101000110",
"100111001",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"010111000",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"001000011",
"101000100",
"101000101",
"100111010",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"001000010",
"101000011",
"101000100",
"100111011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"010111010",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"001000001",
"101000010",
"101000011",
"100111100",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"001000000",
"101000001",
"101000010",
"100111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"010111100",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"000111111",
"101000000",
"101000001",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"000111110",
"100111111",
"101000000",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"010111110",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"000111101",
"100111110",
"100111111",
"101000000",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"000111100",
"100111101",
"100111110",
"101000001",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"011000000",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"000111011",
"100111100",
"100111101",
"101000010",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"000111010",
"100111011",
"100111100",
"101000011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"011000010",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"000111001",
"100111010",
"100111011",
"101000100",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"000111000",
"100111001",
"100111010",
"101000101",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"011000100",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"000110111",
"100111000",
"100111001",
"101000110",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"000110110",
"100110111",
"100111000",
"101000111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"011000110",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"000110101",
"100110110",
"100110111",
"101001000",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"000110100",
"100110101",
"100110110",
"101001001",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"011001000",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"000110011",
"100110100",
"100110101",
"101001010",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"000110010",
"100110011",
"100110100",
"101001011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"011001010",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"000110001",
"100110010",
"100110011",
"101001100",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"000110000",
"100110001",
"100110010",
"101001101",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"011001100",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"000101111",
"100110000",
"100110001",
"101001110",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"000101110",
"100101111",
"100110000",
"101001111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"011001110",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"000101101",
"100101110",
"100101111",
"101010000",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"000101100",
"100101101",
"100101110",
"101010001",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"011010000",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"000101011",
"100101100",
"100101101",
"101010010",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"000101010",
"100101011",
"100101100",
"101010011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"011010010",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"000101001",
"100101010",
"100101011",
"101010100",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"000101000",
"100101001",
"100101010",
"101010101",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"011010100",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"000100111",
"100101000",
"100101001",
"101010110",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"000100110",
"100100111",
"100101000",
"101010111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"011010110",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"000100101",
"100100110",
"100100111",
"101011000",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"000100100",
"100100101",
"100100110",
"101011001",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"011011000",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"000100011",
"100100100",
"100100101",
"101011010",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"000100010",
"100100011",
"100100100",
"101011011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"011011010",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"000100001",
"100100010",
"100100011",
"101011100",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"000100000",
"100100001",
"100100010",
"101011101",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"011011100",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"000011111",
"100100000",
"100100001",
"101011110",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"000011110",
"100011111",
"100100000",
"101011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"011011110",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"000011101",
"100011110",
"100011111",
"101100000",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"000011100",
"100011101",
"100011110",
"101100001",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"011100000",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"000011011",
"100011100",
"100011101",
"101100010",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"000011010",
"100011011",
"100011100",
"101100011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"011100010",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"000011001",
"100011010",
"100011011",
"101100100",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"000011000",
"100011001",
"100011010",
"101100101",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"011100100",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"000010111",
"100011000",
"100011001",
"101100110",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"000010110",
"100010111",
"100011000",
"101100111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"011100110",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"000010101",
"100010110",
"100010111",
"101101000",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"000010100",
"100010101",
"100010110",
"101101001",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"011101000",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"000010011",
"100010100",
"100010101",
"101101010",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"000010010",
"100010011",
"100010100",
"101101011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"011101010",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"000010001",
"100010010",
"100010011",
"101101100",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"000010000",
"100010001",
"100010010",
"101101101",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"011101100",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"000001111",
"100010000",
"100010001",
"101101110",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"000001110",
"100001111",
"100010000",
"101101111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"011101110",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"000001101",
"100001110",
"100001111",
"101110000",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"000001100",
"100001101",
"100001110",
"101110001",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"011110000",
"001110010",
"001110001",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"000001011",
"100001100",
"100001101",
"101110010",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"111110000",
"111110001",
"101110011",
"101110010",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"000001010",
"100001011",
"100001100",
"101110011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"111110000",
"111110001",
"011110010",
"001110100",
"001110011",
"001110010",
"001110001",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"000001001",
"100001010",
"100001011",
"101110100",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"111110000",
"111110001",
"111110010",
"111110011",
"101110101",
"101110100",
"101110011",
"101110010",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"000001000",
"100001001",
"100001010",
"101110101",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"111110000",
"111110001",
"111110010",
"111110011",
"011110100",
"001110110",
"001110101",
"001110100",
"001110011",
"001110010",
"001110001",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"000000111",
"100001000",
"100001001",
"101110110",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"111110000",
"111110001",
"111110010",
"111110011",
"111110100",
"111110101",
"101110111",
"101110110",
"101110101",
"101110100",
"101110011",
"101110010",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"000000110",
"100000111",
"100001000",
"101110111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"111110000",
"111110001",
"111110010",
"111110011",
"111110100",
"111110101",
"011110110",
"001111000",
"001110111",
"001110110",
"001110101",
"001110100",
"001110011",
"001110010",
"001110001",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"000000101",
"100000110",
"100000111",
"101111000",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"111110000",
"111110001",
"111110010",
"111110011",
"111110100",
"111110101",
"111110110",
"111110111",
"101111001",
"101111000",
"101110111",
"101110110",
"101110101",
"101110100",
"101110011",
"101110010",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"000000100",
"100000101",
"100000110",
"101111001",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"111110000",
"111110001",
"111110010",
"111110011",
"111110100",
"111110101",
"111110110",
"111110111",
"011111000",
"001111010",
"001111001",
"001111000",
"001110111",
"001110110",
"001110101",
"001110100",
"001110011",
"001110010",
"001110001",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"000000011",
"100000100",
"100000101",
"101111010",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"111110000",
"111110001",
"111110010",
"111110011",
"111110100",
"111110101",
"111110110",
"111110111",
"111111000",
"111111001",
"101111011",
"101111010",
"101111001",
"101111000",
"101110111",
"101110110",
"101110101",
"101110100",
"101110011",
"101110010",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"000000010",
"100000011",
"100000100",
"101111011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"111110000",
"111110001",
"111110010",
"111110011",
"111110100",
"111110101",
"111110110",
"111110111",
"111111000",
"111111001",
"011111010",
"001111100",
"001111011",
"001111010",
"001111001",
"001111000",
"001110111",
"001110110",
"001110101",
"001110100",
"001110011",
"001110010",
"001110001",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"000000001",
"100000010",
"100000011",
"101111100",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"111110000",
"111110001",
"111110010",
"111110011",
"111110100",
"111110101",
"111110110",
"111110111",
"111111000",
"111111001",
"111111010",
"111111011",
"101111101",
"101111100",
"101111011",
"101111010",
"101111001",
"101111000",
"101110111",
"101110110",
"101110101",
"101110100",
"101110011",
"101110010",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"000000001",
"100000001",
"100000010",
"101111101",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"111110000",
"111110001",
"111110010",
"111110011",
"111110100",
"111110101",
"111110110",
"111110111",
"111111000",
"111111001",
"111111010",
"111111011",
"011111100",
"001111110",
"001111101",
"001111100",
"001111011",
"001111010",
"001111001",
"001111000",
"001110111",
"001110110",
"001110101",
"001110100",
"001110011",
"001110010",
"001110001",
"001110000",
"001101111",
"001101110",
"001101101",
"001101100",
"001101011",
"001101010",
"001101001",
"001101000",
"001100111",
"001100110",
"001100101",
"001100100",
"001100011",
"001100010",
"001100001",
"001100000",
"001011111",
"001011110",
"001011101",
"001011100",
"001011011",
"001011010",
"001011001",
"001011000",
"001010111",
"001010110",
"001010101",
"001010100",
"001010011",
"001010010",
"001010001",
"001010000",
"001001111",
"001001110",
"001001101",
"001001100",
"001001011",
"001001010",
"001001001",
"001001000",
"001000111",
"001000110",
"001000101",
"001000100",
"001000011",
"001000010",
"001000001",
"001000000",
"000111111",
"000111110",
"000111101",
"000111100",
"000111011",
"000111010",
"000111001",
"000111000",
"000110111",
"000110110",
"000110101",
"000110100",
"000110011",
"000110010",
"000110001",
"000110000",
"000101111",
"000101110",
"000101101",
"000101100",
"000101011",
"000101010",
"000101001",
"000101000",
"000100111",
"000100110",
"000100101",
"000100100",
"000100011",
"000100010",
"000100001",
"000100000",
"000011111",
"000011110",
"000011101",
"000011100",
"000011011",
"000011010",
"000011001",
"000011000",
"000010111",
"000010110",
"000010101",
"000010100",
"000010011",
"000010010",
"000010001",
"000010000",
"000001111",
"000001110",
"000001101",
"000001100",
"000001011",
"000001010",
"000001001",
"000001000",
"000000111",
"000000110",
"000000101",
"000000100",
"000000011",
"000000010",
"000000010",
"100000001",
"100000001",
"101111110",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"111110000",
"111110001",
"111110010",
"111110011",
"111110100",
"111110101",
"111110110",
"111110111",
"111111000",
"111111001",
"111111010",
"111111011",
"111111100",
"111111101",
"101111111",
"101111110",
"101111101",
"101111100",
"101111011",
"101111010",
"101111001",
"101111000",
"101110111",
"101110110",
"101110101",
"101110100",
"101110011",
"101110010",
"101110001",
"101110000",
"101101111",
"101101110",
"101101101",
"101101100",
"101101011",
"101101010",
"101101001",
"101101000",
"101100111",
"101100110",
"101100101",
"101100100",
"101100011",
"101100010",
"101100001",
"101100000",
"101011111",
"101011110",
"101011101",
"101011100",
"101011011",
"101011010",
"101011001",
"101011000",
"101010111",
"101010110",
"101010101",
"101010100",
"101010011",
"101010010",
"101010001",
"101010000",
"101001111",
"101001110",
"101001101",
"101001100",
"101001011",
"101001010",
"101001001",
"101001000",
"101000111",
"101000110",
"101000101",
"101000100",
"101000011",
"101000010",
"101000001",
"101000000",
"100111111",
"100111110",
"100111101",
"100111100",
"100111011",
"100111010",
"100111001",
"100111000",
"100110111",
"100110110",
"100110101",
"100110100",
"100110011",
"100110010",
"100110001",
"100110000",
"100101111",
"100101110",
"100101101",
"100101100",
"100101011",
"100101010",
"100101001",
"100101000",
"100100111",
"100100110",
"100100101",
"100100100",
"100100011",
"100100010",
"100100001",
"100100000",
"100011111",
"100011110",
"100011101",
"100011100",
"100011011",
"100011010",
"100011001",
"100011000",
"100010111",
"100010110",
"100010101",
"100010100",
"100010011",
"100010010",
"100010001",
"100010000",
"100001111",
"100001110",
"100001101",
"100001100",
"100001011",
"100001010",
"100001001",
"100001000",
"100000111",
"100000110",
"100000101",
"100000100",
"100000011",
"100000010",
"100000010",
"100000001",
"101111111",
"110000000",
"110000001",
"110000010",
"110000011",
"110000100",
"110000101",
"110000110",
"110000111",
"110001000",
"110001001",
"110001010",
"110001011",
"110001100",
"110001101",
"110001110",
"110001111",
"110010000",
"110010001",
"110010010",
"110010011",
"110010100",
"110010101",
"110010110",
"110010111",
"110011000",
"110011001",
"110011010",
"110011011",
"110011100",
"110011101",
"110011110",
"110011111",
"110100000",
"110100001",
"110100010",
"110100011",
"110100100",
"110100101",
"110100110",
"110100111",
"110101000",
"110101001",
"110101010",
"110101011",
"110101100",
"110101101",
"110101110",
"110101111",
"110110000",
"110110001",
"110110010",
"110110011",
"110110100",
"110110101",
"110110110",
"110110111",
"110111000",
"110111001",
"110111010",
"110111011",
"110111100",
"110111101",
"110111110",
"110111111",
"111000000",
"111000001",
"111000010",
"111000011",
"111000100",
"111000101",
"111000110",
"111000111",
"111001000",
"111001001",
"111001010",
"111001011",
"111001100",
"111001101",
"111001110",
"111001111",
"111010000",
"111010001",
"111010010",
"111010011",
"111010100",
"111010101",
"111010110",
"111010111",
"111011000",
"111011001",
"111011010",
"111011011",
"111011100",
"111011101",
"111011110",
"111011111",
"111100000",
"111100001",
"111100010",
"111100011",
"111100100",
"111100101",
"111100110",
"111100111",
"111101000",
"111101001",
"111101010",
"111101011",
"111101100",
"111101101",
"111101110",
"111101111",
"111110000",
"111110001",
"111110010",
"111110011",
"111110100",
"111110101",
"111110110",
"111110111",
"111111000",
"111111001",
"111111010",
"111111011",
"111111100",
"111111101",
"111111110"
);

begin

    process(clk)
    begin
        if (rising_edge(clk)) then
            sum <= rom(to_integer(unsigned(addr_r)));
        end if;
    end process;

    addr_r <= a & b;
    
end Behavioral;
       
