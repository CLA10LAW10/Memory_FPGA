module fifo
  #(
   parameter DATA_WIDTH=4, // number of bits in a word
             ADDR_WIDTH=4  // number of address bits
  )
  (
   input  logic clk, reset,
   input  logic rd, wr,
   input  logic [DATA_WIDTH-1:0] w_data,
   output logic almost_empty, almost_full,
   output logic empty, full,
   output logic [ADDR_WIDTH+1:0] word_count,
   output logic [DATA_WIDTH-1:0] r_data
  );

  //signal declaration
  logic [ADDR_WIDTH-1:0] w_addr, r_addr;
  logic wr_en, full_tmp;
  // body
  // write enabled only when FIFO is not full
  assign wr_en = wr & ~full_tmp;
  assign full = full_tmp;
 
  // instantiate fifo control unit
  fifo_ctrl #(.ADDR_WIDTH(ADDR_WIDTH)) c_unit
     (.*, .full(full_tmp));

  // instantiate register file
  reg_file
     #(.DATA_WIDTH(DATA_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) f_unit (.*);
endmodule
